----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:11:24 04/10/2016 
-- Design Name: 
-- Module Name:    shift_module - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity shift_module is
    Port ( operand_a : in  STD_LOGIC_VECTOR (15 downto 0);
           operand_b : in  STD_LOGIC_VECTOR (15 downto 0);
			  shamt		: in 	STD_LOGIC_VECTOR(4 downto 0);
           operation : in  STD_LOGIC;
           result 	: out STD_LOGIC_VECTOR (15 downto 0));
end shift_module;

architecture Behavioral of shift_module is

begin
	result <= 	to_stdlogicvector(to_bitvector(operand_a) sll to_integer(unsigned(shamt))) when operation= '0'
		else 		to_stdlogicvector(to_bitvector(operand_a) sll to_integer(unsigned(shamt)));

end Behavioral;

